-------------------------------------------------------------------------------
-- Title      : AES testbench
-- Project    : Extensible Rijndael Block Cipher using VHDL-2008
-------------------------------------------------------------------------------
-- File       : AES_tb.vhd
-- Author     : Clyde R. Visser  <Clyde.R.Visser@gmail.com>
-- Company    : eXpertroniX
-- Created    : 2023-04-23
-- Last update: 2023-04-29
-- Platform   : Modelsim
-- Standard   : VHDL'08, Math Packages
-------------------------------------------------------------------------------
-- Description: AES testbench for ECB, CBC, CFB128, OFB, CTR Modes of Operation
-- using 256, 192, & 128 bit key sizes
-------------------------------------------------------------------------------
--
-- Copyright 2023 eXpertroniX
-- SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
--
-- Licensed under the Solderpad Hardware License v 2.1 (the “License”); you may
-- not use this file except in compliance with the License, or, at your option,
-- the Apache License version 2.0. You may obtain a copy of the License at
-- https://solderpad.org/licenses/SHL-2.1/
--
-- Unless required by applicable law or agreed to in writing, any work
-- distributed under the License is distributed on an “AS IS” BASIS, WITHOUT
-- WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. See the
-- License for the specific language governing permissions and limitations
-- under the License.
--
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2023-04-23  1.0      Clyde   Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.Rijndael.all;
use work.testbench_utils.all;

entity testbench is
end entity testbench;

architecture behavior of testbench is

  constant WordSize  : natural  := 8;
  constant WordRange : natural  := 2**WordSize;
  subtype WordType is FiniteField(WordSize-1 downto 0);
  constant Word      : WordType := (others => '0');

  -----------------------------------------------------------------------------
  -- Test vectors taken from:
  -- NIST Special Publication 800-38A Recommendation for Block 2001 Edition
  -- Cipher Modes of Operation, Methods and Techniques
  -- Appendix F: Example Vectors for Modes of Operation of the AES
  -----------------------------------------------------------------------------

  -- Key: 603deb1015ca71be2b73aef0857d77811f352c073b6108d72d9810a30914dff4
  constant Key256 : KeyType(0 to 8-1)(0 to 4-1)(7 downto 0) := (
    0 => (0 => x"60", 1 => x"3d", 2 => x"eb", 3 => x"10"),  -- 603deb10
    1 => (0 => x"15", 1 => x"ca", 2 => x"71", 3 => x"be"),  -- 15ca71be
    2 => (0 => x"2b", 1 => x"73", 2 => x"ae", 3 => x"f0"),  -- 2b73aef0
    3 => (0 => x"85", 1 => x"7d", 2 => x"77", 3 => x"81"),  -- 857d7781
    4 => (0 => x"1f", 1 => x"35", 2 => x"2c", 3 => x"07"),  -- 1f352c07
    5 => (0 => x"3b", 1 => x"61", 2 => x"08", 3 => x"d7"),  -- 3b6108d7
    6 => (0 => x"2d", 1 => x"98", 2 => x"10", 3 => x"a3"),  -- 2d9810a3
    7 => (0 => x"09", 1 => x"14", 2 => x"df", 3 => x"f4")   -- 0914dff4
    );

  -- Key: 8e73b0f7da0e6452c810f32b809079e562f8ead2522c6b7b
  constant Key192 : KeyType(0 to 6-1)(0 to 4-1)(7 downto 0) := (
    0 => (0 => x"8e", 1 => x"73", 2 => x"b0", 3 => x"f7"),  -- 8e73b0f7
    1 => (0 => x"da", 1 => x"0e", 2 => x"64", 3 => x"52"),  -- da0e6452
    2 => (0 => x"c8", 1 => x"10", 2 => x"f3", 3 => x"2b"),  -- c810f32b
    3 => (0 => x"80", 1 => x"90", 2 => x"79", 3 => x"e5"),  -- 809079e5
    4 => (0 => x"62", 1 => x"f8", 2 => x"ea", 3 => x"d2"),  -- 62f8ead2
    5 => (0 => x"52", 1 => x"2c", 2 => x"6b", 3 => x"7b")   -- 522c6b7b
    );

  -- Key: 2b7e151628aed2a6abf7158809cf4f3c
  constant Key128 : KeyType(0 to 4-1)(0 to 4-1)(7 downto 0) := (
    0 => (0 => x"2b", 1 => x"7e", 2 => x"15", 3 => x"16"),  -- 2b7e1516
    1 => (0 => x"28", 1 => x"ae", 2 => x"d2", 3 => x"a6"),  -- 28aed2a6
    2 => (0 => x"ab", 1 => x"f7", 2 => x"15", 3 => x"88"),  -- abf71588
    3 => (0 => x"09", 1 => x"cf", 2 => x"4f", 3 => x"3c")   -- 09cf4f3c
    );

  -- IV: 000102030405060708090a0b0c0d0e0f
  constant InitializationVector : StateType(0 to 4-1)(0 to 4-1)(7 downto 0) := (
    0 => (0 => x"00", 1 => x"01", 2 => x"02", 3 => x"03"),  -- 00010203
    1 => (0 => x"04", 1 => x"05", 2 => x"06", 3 => x"07"),  -- 04050607
    2 => (0 => x"08", 1 => x"09", 2 => x"0a", 3 => x"0b"),  -- 08090a0b
    3 => (0 => x"0c", 1 => x"0d", 2 => x"0e", 3 => x"0f")   -- 0c0d0e0f
    );

  -- Ctr: f0f1f2f3f4f5f6f7f8f9fafbfcfdfeff
  constant InitialCounter : StateType(0 to 4-1)(0 to 4-1)(7 downto 0) := (
    0 => (0 => x"f0", 1 => x"f1", 2 => x"f2", 3 => x"f3"),  -- f0f1f2f3
    1 => (0 => x"f4", 1 => x"f5", 2 => x"f6", 3 => x"f7"),  -- f4f5f6f7
    2 => (0 => x"f8", 1 => x"f9", 2 => x"fa", 3 => x"fb"),  -- f8f9fafb
    3 => (0 => x"fc", 1 => x"fd", 2 => x"fe", 3 => x"ff")   -- fcfdfeff
    );

  type TestVectorType is array (natural range <>, natural range <>) of StateType;

  constant TestVector256_ECB : TestVectorType(0 to 3, 0 to 1)(0 to 4-1)(0 to 4-1)(7 downto 0) :=
    (
      0 =>
      (
        0 =>
        -- 6bc1bee22e409f96e93d7e117393172a
        (0 => (0 => x"6b", 1 => x"c1", 2 => x"be", 3 => x"e2"),   -- 6bc1bee2
         1 => (0 => x"2e", 1 => x"40", 2 => x"9f", 3 => x"96"),   -- 2e409f96
         2 => (0 => x"e9", 1 => x"3d", 2 => x"7e", 3 => x"11"),   -- e93d7e11
         3 => (0 => x"73", 1 => x"93", 2 => x"17", 3 => x"2a")),  -- 7393172a
        1 =>
        -- f3eed1bdb5d2a03c064b5a7e3db181f8
        (0 => (0 => x"f3", 1 => x"ee", 2 => x"d1", 3 => x"bd"),   -- f3eed1bd
         1 => (0 => x"b5", 1 => x"d2", 2 => x"a0", 3 => x"3c"),   -- b5d2a03c
         2 => (0 => x"06", 1 => x"4b", 2 => x"5a", 3 => x"7e"),   -- 064b5a7e
         3 => (0 => x"3d", 1 => x"b1", 2 => x"81", 3 => x"f8"))   -- 3db181f8
        ),
      1 =>
      (
        0 =>
        -- ae2d8a571e03ac9c9eb76fac45af8e51
        (0 => (0 => x"ae", 1 => x"2d", 2 => x"8a", 3 => x"57"),   -- ae2d8a57
         1 => (0 => x"1e", 1 => x"03", 2 => x"ac", 3 => x"9c"),   -- 1e03ac9c
         2 => (0 => x"9e", 1 => x"b7", 2 => x"6f", 3 => x"ac"),   -- 9eb76fac
         3 => (0 => x"45", 1 => x"af", 2 => x"8e", 3 => x"51")),  -- 45af8e51
        1 =>
        -- 591ccb10d410ed26dc5ba74a31362870
        (0 => (0 => x"59", 1 => x"1c", 2 => x"cb", 3 => x"10"),   -- 591ccb10
         1 => (0 => x"d4", 1 => x"10", 2 => x"ed", 3 => x"26"),   -- d410ed26
         2 => (0 => x"dc", 1 => x"5b", 2 => x"a7", 3 => x"4a"),   -- dc5ba74a
         3 => (0 => x"31", 1 => x"36", 2 => x"28", 3 => x"70"))   -- 31362870
        ),
      2 =>
      (
        0 =>
        -- 30c81c46a35ce411e5fbc1191a0a52ef
        (0 => (0 => x"30", 1 => x"c8", 2 => x"1c", 3 => x"46"),   -- 30c81c46
         1 => (0 => x"a3", 1 => x"5c", 2 => x"e4", 3 => x"11"),   -- a35ce411
         2 => (0 => x"e5", 1 => x"fb", 2 => x"c1", 3 => x"19"),   -- e5fbc119
         3 => (0 => x"1a", 1 => x"0a", 2 => x"52", 3 => x"ef")),  -- 1a0a52ef
        1 =>
        -- b6ed21b99ca6f4f9f153e7b1beafed1d
        (0 => (0 => x"b6", 1 => x"ed", 2 => x"21", 3 => x"b9"),   -- b6ed21b9
         1 => (0 => x"9c", 1 => x"a6", 2 => x"f4", 3 => x"f9"),   -- 9ca6f4f9
         2 => (0 => x"f1", 1 => x"53", 2 => x"e7", 3 => x"b1"),   -- f153e7b1
         3 => (0 => x"be", 1 => x"af", 2 => x"ed", 3 => x"1d"))   -- beafed1d
        ),
      3 =>
      (
        0 =>
        -- f69f2445df4f9b17ad2b417be66c3710
        (0 => (0 => x"f6", 1 => x"9f", 2 => x"24", 3 => x"45"),   -- f69f2445
         1 => (0 => x"df", 1 => x"4f", 2 => x"9b", 3 => x"17"),   -- df4f9b17
         2 => (0 => x"ad", 1 => x"2b", 2 => x"41", 3 => x"7b"),   -- ad2b417b
         3 => (0 => x"e6", 1 => x"6c", 2 => x"37", 3 => x"10")),  -- e66c3710
        1 =>
        -- 23304b7a39f9f3ff067d8d8f9e24ecc7
        (0 => (0 => x"23", 1 => x"30", 2 => x"4b", 3 => x"7a"),   -- 23304b7a
         1 => (0 => x"39", 1 => x"f9", 2 => x"f3", 3 => x"ff"),   -- 39f9f3ff
         2 => (0 => x"06", 1 => x"7d", 2 => x"8d", 3 => x"8f"),   -- 067d8d8f
         3 => (0 => x"9e", 1 => x"24", 2 => x"ec", 3 => x"c7"))   -- 9e24ecc7
        )
      );


  constant TestVector256_CBC : TestVectorType(0 to 3, 0 to 1)(0 to 4-1)(0 to 4-1)(7 downto 0) :=
    (
      0 =>
      (
        0 =>
        -- 6bc1bee22e409f96e93d7e117393172a
        (0 => (0 => x"6b", 1 => x"c1", 2 => x"be", 3 => x"e2"),   -- 6bc1bee2
         1 => (0 => x"2e", 1 => x"40", 2 => x"9f", 3 => x"96"),   -- 2e409f96
         2 => (0 => x"e9", 1 => x"3d", 2 => x"7e", 3 => x"11"),   -- e93d7e11
         3 => (0 => x"73", 1 => x"93", 2 => x"17", 3 => x"2a")),  -- 7393172a
        1 =>
        -- f58c4c04d6e5f1ba779eabfb5f7bfbd6
        (0 => (0 => x"f5", 1 => x"8c", 2 => x"4c", 3 => x"04"),   -- f58c4c04
         1 => (0 => x"d6", 1 => x"e5", 2 => x"f1", 3 => x"ba"),   -- d6e5f1ba
         2 => (0 => x"77", 1 => x"9e", 2 => x"ab", 3 => x"fb"),   -- 779eabfb
         3 => (0 => x"5f", 1 => x"7b", 2 => x"fb", 3 => x"d6"))   -- 5f7bfbd6
        ),
      1 =>
      (
        0 =>
        -- ae2d8a571e03ac9c9eb76fac45af8e51
        (0 => (0 => x"ae", 1 => x"2d", 2 => x"8a", 3 => x"57"),   -- ae2d8a57
         1 => (0 => x"1e", 1 => x"03", 2 => x"ac", 3 => x"9c"),   -- 1e03ac9c
         2 => (0 => x"9e", 1 => x"b7", 2 => x"6f", 3 => x"ac"),   -- 9eb76fac
         3 => (0 => x"45", 1 => x"af", 2 => x"8e", 3 => x"51")),  -- 45af8e51
        1 =>
        -- 9cfc4e967edb808d679f777bc6702c7d
        (0 => (0 => x"9c", 1 => x"fc", 2 => x"4e", 3 => x"96"),   -- 9cfc4e96
         1 => (0 => x"7e", 1 => x"db", 2 => x"80", 3 => x"8d"),   -- 7edb808d
         2 => (0 => x"67", 1 => x"9f", 2 => x"77", 3 => x"7b"),   -- 679f777b
         3 => (0 => x"c6", 1 => x"70", 2 => x"2c", 3 => x"7d"))   -- c6702c7d
        ),
      2 =>
      (
        0 =>
        -- 30c81c46a35ce411e5fbc1191a0a52ef
        (0 => (0 => x"30", 1 => x"c8", 2 => x"1c", 3 => x"46"),   -- 30c81c46
         1 => (0 => x"a3", 1 => x"5c", 2 => x"e4", 3 => x"11"),   -- a35ce411
         2 => (0 => x"e5", 1 => x"fb", 2 => x"c1", 3 => x"19"),   -- e5fbc119
         3 => (0 => x"1a", 1 => x"0a", 2 => x"52", 3 => x"ef")),  -- 1a0a52ef
        1 =>
        -- 39f23369a9d9bacfa530e26304231461
        (0 => (0 => x"39", 1 => x"f2", 2 => x"33", 3 => x"69"),   -- 39f23369
         1 => (0 => x"a9", 1 => x"d9", 2 => x"ba", 3 => x"cf"),   -- a9d9bacf
         2 => (0 => x"a5", 1 => x"30", 2 => x"e2", 3 => x"63"),   -- a530e263
         3 => (0 => x"04", 1 => x"23", 2 => x"14", 3 => x"61"))   -- 04231461
        ),
      3 =>
      (
        0 =>
        -- f69f2445df4f9b17ad2b417be66c3710
        (0 => (0 => x"f6", 1 => x"9f", 2 => x"24", 3 => x"45"),   -- f69f2445
         1 => (0 => x"df", 1 => x"4f", 2 => x"9b", 3 => x"17"),   -- df4f9b17
         2 => (0 => x"ad", 1 => x"2b", 2 => x"41", 3 => x"7b"),   -- ad2b417b
         3 => (0 => x"e6", 1 => x"6c", 2 => x"37", 3 => x"10")),  -- e66c3710
        1 =>
        -- b2eb05e2c39be9fcda6c19078c6a9d1b
        (0 => (0 => x"b2", 1 => x"eb", 2 => x"05", 3 => x"e2"),   -- b2eb05e2
         1 => (0 => x"c3", 1 => x"9b", 2 => x"e9", 3 => x"fc"),   -- c39be9fc
         2 => (0 => x"da", 1 => x"6c", 2 => x"19", 3 => x"07"),   -- da6c1907
         3 => (0 => x"8c", 1 => x"6a", 2 => x"9d", 3 => x"1b"))   -- 8c6a9d1b
        )
      );


  constant TestVector256_CFB128 : TestVectorType(0 to 3, 0 to 1)(0 to 4-1)(0 to 4-1)(7 downto 0) :=
    (
      0 =>
      (
        0 =>
        -- 6bc1bee22e409f96e93d7e117393172a
        (0 => (0 => x"6b", 1 => x"c1", 2 => x"be", 3 => x"e2"),   -- 6bc1bee2
         1 => (0 => x"2e", 1 => x"40", 2 => x"9f", 3 => x"96"),   -- 2e409f96
         2 => (0 => x"e9", 1 => x"3d", 2 => x"7e", 3 => x"11"),   -- e93d7e11
         3 => (0 => x"73", 1 => x"93", 2 => x"17", 3 => x"2a")),  -- 7393172a
        1 =>
        -- dc7e84bfda79164b7ecd8486985d3860
        (0 => (0 => x"dc", 1 => x"7e", 2 => x"84", 3 => x"bf"),   -- dc7e84bf
         1 => (0 => x"da", 1 => x"79", 2 => x"16", 3 => x"4b"),   -- da79164b
         2 => (0 => x"7e", 1 => x"cd", 2 => x"84", 3 => x"86"),   -- 7ecd8486
         3 => (0 => x"98", 1 => x"5d", 2 => x"38", 3 => x"60"))   -- 985d3860
        ),
      1 =>
      (
        0 =>
        -- ae2d8a571e03ac9c9eb76fac45af8e51
        (0 => (0 => x"ae", 1 => x"2d", 2 => x"8a", 3 => x"57"),   -- ae2d8a57
         1 => (0 => x"1e", 1 => x"03", 2 => x"ac", 3 => x"9c"),   -- 1e03ac9c
         2 => (0 => x"9e", 1 => x"b7", 2 => x"6f", 3 => x"ac"),   -- 9eb76fac
         3 => (0 => x"45", 1 => x"af", 2 => x"8e", 3 => x"51")),  -- 45af8e51
        1 =>
        -- 39ffed143b28b1c832113c6331e5407b
        (0 => (0 => x"39", 1 => x"ff", 2 => x"ed", 3 => x"14"),   -- 39ffed14
         1 => (0 => x"3b", 1 => x"28", 2 => x"b1", 3 => x"c8"),   -- 3b28b1c8
         2 => (0 => x"32", 1 => x"11", 2 => x"3c", 3 => x"63"),   -- 32113c63
         3 => (0 => x"31", 1 => x"e5", 2 => x"40", 3 => x"7b"))   -- 31e5407b
        ),
      2 =>
      (
        0 =>
        -- 30c81c46a35ce411e5fbc1191a0a52ef
        (0 => (0 => x"30", 1 => x"c8", 2 => x"1c", 3 => x"46"),   -- 30c81c46
         1 => (0 => x"a3", 1 => x"5c", 2 => x"e4", 3 => x"11"),   -- a35ce411
         2 => (0 => x"e5", 1 => x"fb", 2 => x"c1", 3 => x"19"),   -- e5fbc119
         3 => (0 => x"1a", 1 => x"0a", 2 => x"52", 3 => x"ef")),  -- 1a0a52ef
        1 =>
        -- df10132415e54b92a13ed0a8267ae2f9
        (0 => (0 => x"df", 1 => x"10", 2 => x"13", 3 => x"24"),   -- df101324
         1 => (0 => x"15", 1 => x"e5", 2 => x"4b", 3 => x"92"),   -- 15e54b92
         2 => (0 => x"a1", 1 => x"3e", 2 => x"d0", 3 => x"a8"),   -- a13ed0a8
         3 => (0 => x"26", 1 => x"7a", 2 => x"e2", 3 => x"f9"))   -- 267ae2f9
        ),
      3 =>
      (
        0 =>
        -- f69f2445df4f9b17ad2b417be66c3710
        (0 => (0 => x"f6", 1 => x"9f", 2 => x"24", 3 => x"45"),   -- f69f2445
         1 => (0 => x"df", 1 => x"4f", 2 => x"9b", 3 => x"17"),   -- df4f9b17
         2 => (0 => x"ad", 1 => x"2b", 2 => x"41", 3 => x"7b"),   -- ad2b417b
         3 => (0 => x"e6", 1 => x"6c", 2 => x"37", 3 => x"10")),  -- e66c3710
        1 =>
        -- 75a385741ab9cef82031623d55b1e471
        (0 => (0 => x"75", 1 => x"a3", 2 => x"85", 3 => x"74"),   -- 75a38574
         1 => (0 => x"1a", 1 => x"b9", 2 => x"ce", 3 => x"f8"),   -- 1ab9cef8
         2 => (0 => x"20", 1 => x"31", 2 => x"62", 3 => x"3d"),   -- 2031623d
         3 => (0 => x"55", 1 => x"b1", 2 => x"e4", 3 => x"71"))   -- 55b1e471
        )
      );


  constant TestVector256_OFB : TestVectorType(0 to 3, 0 to 1)(0 to 4-1)(0 to 4-1)(7 downto 0) :=
    (
      0 =>
      (
        0 =>
        -- 6bc1bee22e409f96e93d7e117393172a
        (0 => (0 => x"6b", 1 => x"c1", 2 => x"be", 3 => x"e2"),   -- 6bc1bee2
         1 => (0 => x"2e", 1 => x"40", 2 => x"9f", 3 => x"96"),   -- 2e409f96
         2 => (0 => x"e9", 1 => x"3d", 2 => x"7e", 3 => x"11"),   -- e93d7e11
         3 => (0 => x"73", 1 => x"93", 2 => x"17", 3 => x"2a")),  -- 7393172a
        1 =>
        -- dc7e84bfda79164b7ecd8486985d3860
        (0 => (0 => x"dc", 1 => x"7e", 2 => x"84", 3 => x"bf"),   -- dc7e84bf
         1 => (0 => x"da", 1 => x"79", 2 => x"16", 3 => x"4b"),   -- da79164b
         2 => (0 => x"7e", 1 => x"cd", 2 => x"84", 3 => x"86"),   -- 7ecd8486
         3 => (0 => x"98", 1 => x"5d", 2 => x"38", 3 => x"60"))   -- 985d3860
        ),
      1 =>
      (
        0 =>
        -- ae2d8a571e03ac9c9eb76fac45af8e51
        (0 => (0 => x"ae", 1 => x"2d", 2 => x"8a", 3 => x"57"),   -- ae2d8a57
         1 => (0 => x"1e", 1 => x"03", 2 => x"ac", 3 => x"9c"),   -- 1e03ac9c
         2 => (0 => x"9e", 1 => x"b7", 2 => x"6f", 3 => x"ac"),   -- 9eb76fac
         3 => (0 => x"45", 1 => x"af", 2 => x"8e", 3 => x"51")),  -- 45af8e51
        1 =>
        -- 4febdc6740d20b3ac88f6ad82a4fb08d
        (0 => (0 => x"4f", 1 => x"eb", 2 => x"dc", 3 => x"67"),   -- 4febdc67
         1 => (0 => x"40", 1 => x"d2", 2 => x"0b", 3 => x"3a"),   -- 40d20b3a
         2 => (0 => x"c8", 1 => x"8f", 2 => x"6a", 3 => x"d8"),   -- c88f6ad8
         3 => (0 => x"2a", 1 => x"4f", 2 => x"b0", 3 => x"8d"))   -- 2a4fb08d
        ),
      2 =>
      (
        0 =>
        -- 30c81c46a35ce411e5fbc1191a0a52ef
        (0 => (0 => x"30", 1 => x"c8", 2 => x"1c", 3 => x"46"),   -- 30c81c46
         1 => (0 => x"a3", 1 => x"5c", 2 => x"e4", 3 => x"11"),   -- a35ce411
         2 => (0 => x"e5", 1 => x"fb", 2 => x"c1", 3 => x"19"),   -- e5fbc119
         3 => (0 => x"1a", 1 => x"0a", 2 => x"52", 3 => x"ef")),  -- 1a0a52ef
        1 =>
        -- 71ab47a086e86eedf39d1c5bba97c408
        (0 => (0 => x"71", 1 => x"ab", 2 => x"47", 3 => x"a0"),   -- 71ab47a0
         1 => (0 => x"86", 1 => x"e8", 2 => x"6e", 3 => x"ed"),   -- 86e86eed
         2 => (0 => x"f3", 1 => x"9d", 2 => x"1c", 3 => x"5b"),   -- f39d1c5b
         3 => (0 => x"ba", 1 => x"97", 2 => x"c4", 3 => x"08"))   -- ba97c408
        ),
      3 =>
      (
        0 =>
        -- f69f2445df4f9b17ad2b417be66c3710
        (0 => (0 => x"f6", 1 => x"9f", 2 => x"24", 3 => x"45"),   -- f69f2445
         1 => (0 => x"df", 1 => x"4f", 2 => x"9b", 3 => x"17"),   -- df4f9b17
         2 => (0 => x"ad", 1 => x"2b", 2 => x"41", 3 => x"7b"),   -- ad2b417b
         3 => (0 => x"e6", 1 => x"6c", 2 => x"37", 3 => x"10")),  -- e66c3710
        1 =>
        -- 0126141d67f37be8538f5a8be740e484
        (0 => (0 => x"01", 1 => x"26", 2 => x"14", 3 => x"1d"),   -- 0126141d
         1 => (0 => x"67", 1 => x"f3", 2 => x"7b", 3 => x"e8"),   -- 67f37be8
         2 => (0 => x"53", 1 => x"8f", 2 => x"5a", 3 => x"8b"),   -- 538f5a8b
         3 => (0 => x"e7", 1 => x"40", 2 => x"e4", 3 => x"84"))   -- e740e484
        )
      );


  constant TestVector256_CTR : TestVectorType(0 to 3, 0 to 1)(0 to 4-1)(0 to 4-1)(7 downto 0) :=
    (
      0 =>
      (
        0 =>
        -- 6bc1bee22e409f96e93d7e117393172a
        (0 => (0 => x"6b", 1 => x"c1", 2 => x"be", 3 => x"e2"),   -- 6bc1bee2
         1 => (0 => x"2e", 1 => x"40", 2 => x"9f", 3 => x"96"),   -- 2e409f96
         2 => (0 => x"e9", 1 => x"3d", 2 => x"7e", 3 => x"11"),   -- e93d7e11
         3 => (0 => x"73", 1 => x"93", 2 => x"17", 3 => x"2a")),  -- 7393172a
        1 =>
        -- 601ec313775789a5b7a7f504bbf3d228
        (0 => (0 => x"60", 1 => x"1e", 2 => x"c3", 3 => x"13"),   -- 601ec313
         1 => (0 => x"77", 1 => x"57", 2 => x"89", 3 => x"a5"),   -- 775789a5
         2 => (0 => x"b7", 1 => x"a7", 2 => x"f5", 3 => x"04"),   -- b7a7f504
         3 => (0 => x"bb", 1 => x"f3", 2 => x"d2", 3 => x"28"))   -- bbf3d228
        ),
      1 =>
      (
        0 =>
        -- ae2d8a571e03ac9c9eb76fac45af8e51
        (0 => (0 => x"ae", 1 => x"2d", 2 => x"8a", 3 => x"57"),   -- ae2d8a57
         1 => (0 => x"1e", 1 => x"03", 2 => x"ac", 3 => x"9c"),   -- 1e03ac9c
         2 => (0 => x"9e", 1 => x"b7", 2 => x"6f", 3 => x"ac"),   -- 9eb76fac
         3 => (0 => x"45", 1 => x"af", 2 => x"8e", 3 => x"51")),  -- 45af8e51
        1 =>
        -- f443e3ca4d62b59aca84e990cacaf5c5
        (0 => (0 => x"f4", 1 => x"43", 2 => x"e3", 3 => x"ca"),   -- f443e3ca
         1 => (0 => x"4d", 1 => x"62", 2 => x"b5", 3 => x"9a"),   -- 4d62b59a
         2 => (0 => x"ca", 1 => x"84", 2 => x"e9", 3 => x"90"),   -- ca84e990
         3 => (0 => x"ca", 1 => x"ca", 2 => x"f5", 3 => x"c5"))   -- cacaf5c5
        ),
      2 =>
      (
        0 =>
        -- 30c81c46a35ce411e5fbc1191a0a52ef
        (0 => (0 => x"30", 1 => x"c8", 2 => x"1c", 3 => x"46"),   -- 30c81c46
         1 => (0 => x"a3", 1 => x"5c", 2 => x"e4", 3 => x"11"),   -- a35ce411
         2 => (0 => x"e5", 1 => x"fb", 2 => x"c1", 3 => x"19"),   -- e5fbc119
         3 => (0 => x"1a", 1 => x"0a", 2 => x"52", 3 => x"ef")),  -- 1a0a52ef
        1 =>
        -- 2b0930daa23de94ce87017ba2d84988d
        (0 => (0 => x"2b", 1 => x"09", 2 => x"30", 3 => x"da"),   -- 2b0930da
         1 => (0 => x"a2", 1 => x"3d", 2 => x"e9", 3 => x"4c"),   -- a23de94c
         2 => (0 => x"e8", 1 => x"70", 2 => x"17", 3 => x"ba"),   -- e87017ba
         3 => (0 => x"2d", 1 => x"84", 2 => x"98", 3 => x"8d"))   -- 2d84988d
        ),
      3 =>
      (
        0 =>
        -- f69f2445df4f9b17ad2b417be66c3710
        (0 => (0 => x"f6", 1 => x"9f", 2 => x"24", 3 => x"45"),   -- f69f2445
         1 => (0 => x"df", 1 => x"4f", 2 => x"9b", 3 => x"17"),   -- df4f9b17
         2 => (0 => x"ad", 1 => x"2b", 2 => x"41", 3 => x"7b"),   -- ad2b417b
         3 => (0 => x"e6", 1 => x"6c", 2 => x"37", 3 => x"10")),  -- e66c3710
        1 =>
        -- dfc9c58db67aada613c2dd08457941a6
        (0 => (0 => x"df", 1 => x"c9", 2 => x"c5", 3 => x"8d"),   -- dfc9c58d
         1 => (0 => x"b6", 1 => x"7a", 2 => x"ad", 3 => x"a6"),   -- b67aada6
         2 => (0 => x"13", 1 => x"c2", 2 => x"dd", 3 => x"08"),   -- 13c2dd08
         3 => (0 => x"45", 1 => x"79", 2 => x"41", 3 => x"a6"))   -- 457941a6
        )
      );


  constant TestVector192_ECB : TestVectorType(0 to 3, 0 to 1)(0 to 4-1)(0 to 4-1)(7 downto 0) :=
    (
      0 =>
      (
        0 =>
        -- 6bc1bee22e409f96e93d7e117393172a
        (0 => (0 => x"6b", 1 => x"c1", 2 => x"be", 3 => x"e2"),   -- 6bc1bee2
         1 => (0 => x"2e", 1 => x"40", 2 => x"9f", 3 => x"96"),   -- 2e409f96
         2 => (0 => x"e9", 1 => x"3d", 2 => x"7e", 3 => x"11"),   -- e93d7e11
         3 => (0 => x"73", 1 => x"93", 2 => x"17", 3 => x"2a")),  -- 7393172a
        1 =>
        -- bd334f1d6e45f25ff712a214571fa5cc
        (0 => (0 => x"bd", 1 => x"33", 2 => x"4f", 3 => x"1d"),   -- bd334f1d
         1 => (0 => x"6e", 1 => x"45", 2 => x"f2", 3 => x"5f"),   -- 6e45f25f
         2 => (0 => x"f7", 1 => x"12", 2 => x"a2", 3 => x"14"),   -- f712a214
         3 => (0 => x"57", 1 => x"1f", 2 => x"a5", 3 => x"cc"))   -- 571fa5cc
        ),
      1 =>
      (
        0 =>
        -- ae2d8a571e03ac9c9eb76fac45af8e51
        (0 => (0 => x"ae", 1 => x"2d", 2 => x"8a", 3 => x"57"),   -- ae2d8a57
         1 => (0 => x"1e", 1 => x"03", 2 => x"ac", 3 => x"9c"),   -- 1e03ac9c
         2 => (0 => x"9e", 1 => x"b7", 2 => x"6f", 3 => x"ac"),   -- 9eb76fac
         3 => (0 => x"45", 1 => x"af", 2 => x"8e", 3 => x"51")),  -- 45af8e51
        1 =>
        -- 974104846d0ad3ad7734ecb3ecee4eef
        (0 => (0 => x"97", 1 => x"41", 2 => x"04", 3 => x"84"),   -- 97410484
         1 => (0 => x"6d", 1 => x"0a", 2 => x"d3", 3 => x"ad"),   -- 6d0ad3ad
         2 => (0 => x"77", 1 => x"34", 2 => x"ec", 3 => x"b3"),   -- 7734ecb3
         3 => (0 => x"ec", 1 => x"ee", 2 => x"4e", 3 => x"ef"))   -- ecee4eef
        ),
      2 =>
      (
        0 =>
        -- 30c81c46a35ce411e5fbc1191a0a52ef
        (0 => (0 => x"30", 1 => x"c8", 2 => x"1c", 3 => x"46"),   -- 30c81c46
         1 => (0 => x"a3", 1 => x"5c", 2 => x"e4", 3 => x"11"),   -- a35ce411
         2 => (0 => x"e5", 1 => x"fb", 2 => x"c1", 3 => x"19"),   -- e5fbc119
         3 => (0 => x"1a", 1 => x"0a", 2 => x"52", 3 => x"ef")),  -- 1a0a52ef
        1 =>
        -- ef7afd2270e2e60adce0ba2face6444e
        (0 => (0 => x"ef", 1 => x"7a", 2 => x"fd", 3 => x"22"),   -- ef7afd22
         1 => (0 => x"70", 1 => x"e2", 2 => x"e6", 3 => x"0a"),   -- 70e2e60a
         2 => (0 => x"dc", 1 => x"e0", 2 => x"ba", 3 => x"2f"),   -- dce0ba2f
         3 => (0 => x"ac", 1 => x"e6", 2 => x"44", 3 => x"4e"))   -- ace6444e
        ),
      3 =>
      (
        0 =>
        -- f69f2445df4f9b17ad2b417be66c3710
        (0 => (0 => x"f6", 1 => x"9f", 2 => x"24", 3 => x"45"),   -- f69f2445
         1 => (0 => x"df", 1 => x"4f", 2 => x"9b", 3 => x"17"),   -- df4f9b17
         2 => (0 => x"ad", 1 => x"2b", 2 => x"41", 3 => x"7b"),   -- ad2b417b
         3 => (0 => x"e6", 1 => x"6c", 2 => x"37", 3 => x"10")),  -- e66c3710
        1 =>
        -- 9a4b41ba738d6c72fb16691603c18e0e
        (0 => (0 => x"9a", 1 => x"4b", 2 => x"41", 3 => x"ba"),   -- 9a4b41ba
         1 => (0 => x"73", 1 => x"8d", 2 => x"6c", 3 => x"72"),   -- 738d6c72
         2 => (0 => x"fb", 1 => x"16", 2 => x"69", 3 => x"16"),   -- fb166916
         3 => (0 => x"03", 1 => x"c1", 2 => x"8e", 3 => x"0e"))   -- 03c18e0e
        )
      );


  constant TestVector192_CBC : TestVectorType(0 to 3, 0 to 1)(0 to 4-1)(0 to 4-1)(7 downto 0) :=
    (
      0 =>
      (
        0 =>
        -- 6bc1bee22e409f96e93d7e117393172a
        (0 => (0 => x"6b", 1 => x"c1", 2 => x"be", 3 => x"e2"),   -- 6bc1bee2
         1 => (0 => x"2e", 1 => x"40", 2 => x"9f", 3 => x"96"),   -- 2e409f96
         2 => (0 => x"e9", 1 => x"3d", 2 => x"7e", 3 => x"11"),   -- e93d7e11
         3 => (0 => x"73", 1 => x"93", 2 => x"17", 3 => x"2a")),  -- 7393172a
        1 =>
        -- 4f021db243bc633d7178183a9fa071e8
        (0 => (0 => x"4f", 1 => x"02", 2 => x"1d", 3 => x"b2"),   -- 4f021db2
         1 => (0 => x"43", 1 => x"bc", 2 => x"63", 3 => x"3d"),   -- 43bc633d
         2 => (0 => x"71", 1 => x"78", 2 => x"18", 3 => x"3a"),   -- 7178183a
         3 => (0 => x"9f", 1 => x"a0", 2 => x"71", 3 => x"e8"))   -- 9fa071e8
        ),
      1 =>
      (
        0 =>
        -- ae2d8a571e03ac9c9eb76fac45af8e51
        (0 => (0 => x"ae", 1 => x"2d", 2 => x"8a", 3 => x"57"),   -- ae2d8a57
         1 => (0 => x"1e", 1 => x"03", 2 => x"ac", 3 => x"9c"),   -- 1e03ac9c
         2 => (0 => x"9e", 1 => x"b7", 2 => x"6f", 3 => x"ac"),   -- 9eb76fac
         3 => (0 => x"45", 1 => x"af", 2 => x"8e", 3 => x"51")),  -- 45af8e51
        1 =>
        -- b4d9ada9ad7dedf4e5e738763f69145a
        (0 => (0 => x"b4", 1 => x"d9", 2 => x"ad", 3 => x"a9"),   -- b4d9ada9
         1 => (0 => x"ad", 1 => x"7d", 2 => x"ed", 3 => x"f4"),   -- ad7dedf4
         2 => (0 => x"e5", 1 => x"e7", 2 => x"38", 3 => x"76"),   -- e5e73876
         3 => (0 => x"3f", 1 => x"69", 2 => x"14", 3 => x"5a"))   -- 3f69145a
        ),
      2 =>
      (
        0 =>
        -- 30c81c46a35ce411e5fbc1191a0a52ef
        (0 => (0 => x"30", 1 => x"c8", 2 => x"1c", 3 => x"46"),   -- 30c81c46
         1 => (0 => x"a3", 1 => x"5c", 2 => x"e4", 3 => x"11"),   -- a35ce411
         2 => (0 => x"e5", 1 => x"fb", 2 => x"c1", 3 => x"19"),   -- e5fbc119
         3 => (0 => x"1a", 1 => x"0a", 2 => x"52", 3 => x"ef")),  -- 1a0a52ef
        1 =>
        -- 571b242012fb7ae07fa9baac3df102e0
        (0 => (0 => x"57", 1 => x"1b", 2 => x"24", 3 => x"20"),   -- 571b2420
         1 => (0 => x"12", 1 => x"fb", 2 => x"7a", 3 => x"e0"),   -- 12fb7ae0
         2 => (0 => x"7f", 1 => x"a9", 2 => x"ba", 3 => x"ac"),   -- 7fa9baac
         3 => (0 => x"3d", 1 => x"f1", 2 => x"02", 3 => x"e0"))   -- 3df102e0
        ),
      3 =>
      (
        0 =>
        -- f69f2445df4f9b17ad2b417be66c3710
        (0 => (0 => x"f6", 1 => x"9f", 2 => x"24", 3 => x"45"),   -- f69f2445
         1 => (0 => x"df", 1 => x"4f", 2 => x"9b", 3 => x"17"),   -- df4f9b17
         2 => (0 => x"ad", 1 => x"2b", 2 => x"41", 3 => x"7b"),   -- ad2b417b
         3 => (0 => x"e6", 1 => x"6c", 2 => x"37", 3 => x"10")),  -- e66c3710
        1 =>
        -- 08b0e27988598881d920a9e64f5615cd
        (0 => (0 => x"08", 1 => x"b0", 2 => x"e2", 3 => x"79"),   -- 08b0e279
         1 => (0 => x"88", 1 => x"59", 2 => x"88", 3 => x"81"),   -- 88598881
         2 => (0 => x"d9", 1 => x"20", 2 => x"a9", 3 => x"e6"),   -- d920a9e6
         3 => (0 => x"4f", 1 => x"56", 2 => x"15", 3 => x"cd"))   -- 4f5615cd
        )
      );


  constant TestVector192_CFB128 : TestVectorType(0 to 3, 0 to 1)(0 to 4-1)(0 to 4-1)(7 downto 0) :=
    (
      0 =>
      (
        0 =>
        -- 6bc1bee22e409f96e93d7e117393172a
        (0 => (0 => x"6b", 1 => x"c1", 2 => x"be", 3 => x"e2"),   -- 6bc1bee2
         1 => (0 => x"2e", 1 => x"40", 2 => x"9f", 3 => x"96"),   -- 2e409f96
         2 => (0 => x"e9", 1 => x"3d", 2 => x"7e", 3 => x"11"),   -- e93d7e11
         3 => (0 => x"73", 1 => x"93", 2 => x"17", 3 => x"2a")),  -- 7393172a
        1 =>
        -- cdc80d6fddf18cab34c25909c99a4174
        (0 => (0 => x"cd", 1 => x"c8", 2 => x"0d", 3 => x"6f"),   -- cdc80d6f
         1 => (0 => x"dd", 1 => x"f1", 2 => x"8c", 3 => x"ab"),   -- ddf18cab
         2 => (0 => x"34", 1 => x"c2", 2 => x"59", 3 => x"09"),   -- 34c25909
         3 => (0 => x"c9", 1 => x"9a", 2 => x"41", 3 => x"74"))   -- c99a4174
        ),
      1 =>
      (
        0 =>
        -- ae2d8a571e03ac9c9eb76fac45af8e51
        (0 => (0 => x"ae", 1 => x"2d", 2 => x"8a", 3 => x"57"),   -- ae2d8a57
         1 => (0 => x"1e", 1 => x"03", 2 => x"ac", 3 => x"9c"),   -- 1e03ac9c
         2 => (0 => x"9e", 1 => x"b7", 2 => x"6f", 3 => x"ac"),   -- 9eb76fac
         3 => (0 => x"45", 1 => x"af", 2 => x"8e", 3 => x"51")),  -- 45af8e51
        1 =>
        -- 67ce7f7f81173621961a2b70171d3d7a
        (0 => (0 => x"67", 1 => x"ce", 2 => x"7f", 3 => x"7f"),   -- 67ce7f7f
         1 => (0 => x"81", 1 => x"17", 2 => x"36", 3 => x"21"),   -- 81173621
         2 => (0 => x"96", 1 => x"1a", 2 => x"2b", 3 => x"70"),   -- 961a2b70
         3 => (0 => x"17", 1 => x"1d", 2 => x"3d", 3 => x"7a"))   -- 171d3d7a
        ),
      2 =>
      (
        0 =>
        -- 30c81c46a35ce411e5fbc1191a0a52ef
        (0 => (0 => x"30", 1 => x"c8", 2 => x"1c", 3 => x"46"),   -- 30c81c46
         1 => (0 => x"a3", 1 => x"5c", 2 => x"e4", 3 => x"11"),   -- a35ce411
         2 => (0 => x"e5", 1 => x"fb", 2 => x"c1", 3 => x"19"),   -- e5fbc119
         3 => (0 => x"1a", 1 => x"0a", 2 => x"52", 3 => x"ef")),  -- 1a0a52ef
        1 =>
        -- 2e1e8a1dd59b88b1c8e60fed1efac4c9
        (0 => (0 => x"2e", 1 => x"1e", 2 => x"8a", 3 => x"1d"),   -- 2e1e8a1d
         1 => (0 => x"d5", 1 => x"9b", 2 => x"88", 3 => x"b1"),   -- d59b88b1
         2 => (0 => x"c8", 1 => x"e6", 2 => x"0f", 3 => x"ed"),   -- c8e60fed
         3 => (0 => x"1e", 1 => x"fa", 2 => x"c4", 3 => x"c9"))   -- 1efac4c9
        ),
      3 =>
      (
        0 =>
        -- f69f2445df4f9b17ad2b417be66c3710
        (0 => (0 => x"f6", 1 => x"9f", 2 => x"24", 3 => x"45"),   -- f69f2445
         1 => (0 => x"df", 1 => x"4f", 2 => x"9b", 3 => x"17"),   -- df4f9b17
         2 => (0 => x"ad", 1 => x"2b", 2 => x"41", 3 => x"7b"),   -- ad2b417b
         3 => (0 => x"e6", 1 => x"6c", 2 => x"37", 3 => x"10")),  -- e66c3710
        1 =>
        -- c05f9f9ca9834fa042ae8fba584b09ff
        (0 => (0 => x"c0", 1 => x"5f", 2 => x"9f", 3 => x"9c"),   -- c05f9f9c
         1 => (0 => x"a9", 1 => x"83", 2 => x"4f", 3 => x"a0"),   -- a9834fa0
         2 => (0 => x"42", 1 => x"ae", 2 => x"8f", 3 => x"ba"),   -- 42ae8fba
         3 => (0 => x"58", 1 => x"4b", 2 => x"09", 3 => x"ff"))   -- 584b09ff
        )
      );


  constant TestVector192_OFB : TestVectorType(0 to 3, 0 to 1)(0 to 4-1)(0 to 4-1)(7 downto 0) :=
    (
      0 =>
      (
        0 =>
        -- 6bc1bee22e409f96e93d7e117393172a
        (0 => (0 => x"6b", 1 => x"c1", 2 => x"be", 3 => x"e2"),   -- 6bc1bee2
         1 => (0 => x"2e", 1 => x"40", 2 => x"9f", 3 => x"96"),   -- 2e409f96
         2 => (0 => x"e9", 1 => x"3d", 2 => x"7e", 3 => x"11"),   -- e93d7e11
         3 => (0 => x"73", 1 => x"93", 2 => x"17", 3 => x"2a")),  -- 7393172a
        1 =>
        -- cdc80d6fddf18cab34c25909c99a4174
        (0 => (0 => x"cd", 1 => x"c8", 2 => x"0d", 3 => x"6f"),   -- cdc80d6f
         1 => (0 => x"dd", 1 => x"f1", 2 => x"8c", 3 => x"ab"),   -- ddf18cab
         2 => (0 => x"34", 1 => x"c2", 2 => x"59", 3 => x"09"),   -- 34c25909
         3 => (0 => x"c9", 1 => x"9a", 2 => x"41", 3 => x"74"))   -- c99a4174
        ),
      1 =>
      (
        0 =>
        -- ae2d8a571e03ac9c9eb76fac45af8e51
        (0 => (0 => x"ae", 1 => x"2d", 2 => x"8a", 3 => x"57"),   -- ae2d8a57
         1 => (0 => x"1e", 1 => x"03", 2 => x"ac", 3 => x"9c"),   -- 1e03ac9c
         2 => (0 => x"9e", 1 => x"b7", 2 => x"6f", 3 => x"ac"),   -- 9eb76fac
         3 => (0 => x"45", 1 => x"af", 2 => x"8e", 3 => x"51")),  -- 45af8e51
        1 =>
        -- fcc28b8d4c63837c09e81700c1100401
        (0 => (0 => x"fc", 1 => x"c2", 2 => x"8b", 3 => x"8d"),   -- fcc28b8d
         1 => (0 => x"4c", 1 => x"63", 2 => x"83", 3 => x"7c"),   -- 4c63837c
         2 => (0 => x"09", 1 => x"e8", 2 => x"17", 3 => x"00"),   -- 09e81700
         3 => (0 => x"c1", 1 => x"10", 2 => x"04", 3 => x"01"))   -- c1100401
        ),
      2 =>
      (
        0 =>
        -- 30c81c46a35ce411e5fbc1191a0a52ef
        (0 => (0 => x"30", 1 => x"c8", 2 => x"1c", 3 => x"46"),   -- 30c81c46
         1 => (0 => x"a3", 1 => x"5c", 2 => x"e4", 3 => x"11"),   -- a35ce411
         2 => (0 => x"e5", 1 => x"fb", 2 => x"c1", 3 => x"19"),   -- e5fbc119
         3 => (0 => x"1a", 1 => x"0a", 2 => x"52", 3 => x"ef")),  -- 1a0a52ef
        1 =>
        -- 8d9a9aeac0f6596f559c6d4daf59a5f2
        (0 => (0 => x"8d", 1 => x"9a", 2 => x"9a", 3 => x"ea"),   -- 8d9a9aea
         1 => (0 => x"c0", 1 => x"f6", 2 => x"59", 3 => x"6f"),   -- c0f6596f
         2 => (0 => x"55", 1 => x"9c", 2 => x"6d", 3 => x"4d"),   -- 559c6d4d
         3 => (0 => x"af", 1 => x"59", 2 => x"a5", 3 => x"f2"))   -- af59a5f2
        ),
      3 =>
      (
        0 =>
        -- f69f2445df4f9b17ad2b417be66c3710
        (0 => (0 => x"f6", 1 => x"9f", 2 => x"24", 3 => x"45"),   -- f69f2445
         1 => (0 => x"df", 1 => x"4f", 2 => x"9b", 3 => x"17"),   -- df4f9b17
         2 => (0 => x"ad", 1 => x"2b", 2 => x"41", 3 => x"7b"),   -- ad2b417b
         3 => (0 => x"e6", 1 => x"6c", 2 => x"37", 3 => x"10")),  -- e66c3710
        1 =>
        -- 6d9f200857ca6c3e9cac524bd9acc92a
        (0 => (0 => x"6d", 1 => x"9f", 2 => x"20", 3 => x"08"),   -- 6d9f2008
         1 => (0 => x"57", 1 => x"ca", 2 => x"6c", 3 => x"3e"),   -- 57ca6c3e
         2 => (0 => x"9c", 1 => x"ac", 2 => x"52", 3 => x"4b"),   -- 9cac524b
         3 => (0 => x"d9", 1 => x"ac", 2 => x"c9", 3 => x"2a"))   -- d9acc92a
        )
      );


  constant TestVector192_CTR : TestVectorType(0 to 3, 0 to 1)(0 to 4-1)(0 to 4-1)(7 downto 0) :=
    (
      0 =>
      (
        0 =>
        -- 6bc1bee22e409f96e93d7e117393172a
        (0 => (0 => x"6b", 1 => x"c1", 2 => x"be", 3 => x"e2"),   -- 6bc1bee2
         1 => (0 => x"2e", 1 => x"40", 2 => x"9f", 3 => x"96"),   -- 2e409f96
         2 => (0 => x"e9", 1 => x"3d", 2 => x"7e", 3 => x"11"),   -- e93d7e11
         3 => (0 => x"73", 1 => x"93", 2 => x"17", 3 => x"2a")),  -- 7393172a
        1 =>
        -- 1abc932417521ca24f2b0459fe7e6e0b
        (0 => (0 => x"1a", 1 => x"bc", 2 => x"93", 3 => x"24"),   -- 1abc9324
         1 => (0 => x"17", 1 => x"52", 2 => x"1c", 3 => x"a2"),   -- 17521ca2
         2 => (0 => x"4f", 1 => x"2b", 2 => x"04", 3 => x"59"),   -- 4f2b0459
         3 => (0 => x"fe", 1 => x"7e", 2 => x"6e", 3 => x"0b"))   -- fe7e6e0b
        ),
      1 =>
      (
        0 =>
        -- ae2d8a571e03ac9c9eb76fac45af8e51
        (0 => (0 => x"ae", 1 => x"2d", 2 => x"8a", 3 => x"57"),   -- ae2d8a57
         1 => (0 => x"1e", 1 => x"03", 2 => x"ac", 3 => x"9c"),   -- 1e03ac9c
         2 => (0 => x"9e", 1 => x"b7", 2 => x"6f", 3 => x"ac"),   -- 9eb76fac
         3 => (0 => x"45", 1 => x"af", 2 => x"8e", 3 => x"51")),  -- 45af8e51
        1 =>
        -- 090339ec0aa6faefd5ccc2c6f4ce8e94
        (0 => (0 => x"09", 1 => x"03", 2 => x"39", 3 => x"ec"),   -- 090339ec
         1 => (0 => x"0a", 1 => x"a6", 2 => x"fa", 3 => x"ef"),   -- 0aa6faef
         2 => (0 => x"d5", 1 => x"cc", 2 => x"c2", 3 => x"c6"),   -- d5ccc2c6
         3 => (0 => x"f4", 1 => x"ce", 2 => x"8e", 3 => x"94"))   -- f4ce8e94
        ),
      2 =>
      (
        0 =>
        -- 30c81c46a35ce411e5fbc1191a0a52ef
        (0 => (0 => x"30", 1 => x"c8", 2 => x"1c", 3 => x"46"),   -- 30c81c46
         1 => (0 => x"a3", 1 => x"5c", 2 => x"e4", 3 => x"11"),   -- a35ce411
         2 => (0 => x"e5", 1 => x"fb", 2 => x"c1", 3 => x"19"),   -- e5fbc119
         3 => (0 => x"1a", 1 => x"0a", 2 => x"52", 3 => x"ef")),  -- 1a0a52ef
        1 =>
        -- 1e36b26bd1ebc670d1bd1d665620abf7
        (0 => (0 => x"1e", 1 => x"36", 2 => x"b2", 3 => x"6b"),   -- 1e36b26b
         1 => (0 => x"d1", 1 => x"eb", 2 => x"c6", 3 => x"70"),   -- d1ebc670
         2 => (0 => x"d1", 1 => x"bd", 2 => x"1d", 3 => x"66"),   -- d1bd1d66
         3 => (0 => x"56", 1 => x"20", 2 => x"ab", 3 => x"f7"))   -- 5620abf7
        ),
      3 =>
      (
        0 =>
        -- f69f2445df4f9b17ad2b417be66c3710
        (0 => (0 => x"f6", 1 => x"9f", 2 => x"24", 3 => x"45"),   -- f69f2445
         1 => (0 => x"df", 1 => x"4f", 2 => x"9b", 3 => x"17"),   -- df4f9b17
         2 => (0 => x"ad", 1 => x"2b", 2 => x"41", 3 => x"7b"),   -- ad2b417b
         3 => (0 => x"e6", 1 => x"6c", 2 => x"37", 3 => x"10")),  -- e66c3710
        1 =>
        -- 4f78a7f6d29809585a97daec58c6b050
        (0 => (0 => x"4f", 1 => x"78", 2 => x"a7", 3 => x"f6"),   -- 4f78a7f6
         1 => (0 => x"d2", 1 => x"98", 2 => x"09", 3 => x"58"),   -- d2980958
         2 => (0 => x"5a", 1 => x"97", 2 => x"da", 3 => x"ec"),   -- 5a97daec
         3 => (0 => x"58", 1 => x"c6", 2 => x"b0", 3 => x"50"))   -- 58c6b050
        )
      );


  constant TestVector128_ECB : TestVectorType(0 to 3, 0 to 1)(0 to 4-1)(0 to 4-1)(7 downto 0) :=
    (
      0 =>
      (
        0 =>
        -- 6bc1bee22e409f96e93d7e117393172a
        (0 => (0 => x"6b", 1 => x"c1", 2 => x"be", 3 => x"e2"),   -- 6bc1bee2
         1 => (0 => x"2e", 1 => x"40", 2 => x"9f", 3 => x"96"),   -- 2e409f96
         2 => (0 => x"e9", 1 => x"3d", 2 => x"7e", 3 => x"11"),   -- e93d7e11
         3 => (0 => x"73", 1 => x"93", 2 => x"17", 3 => x"2a")),  -- 7393172a
        1 =>
        -- 3ad77bb40d7a3660a89ecaf32466ef97
        (0 => (0 => x"3a", 1 => x"d7", 2 => x"7b", 3 => x"b4"),   -- 3ad77bb4
         1 => (0 => x"0d", 1 => x"7a", 2 => x"36", 3 => x"60"),   -- 0d7a3660
         2 => (0 => x"a8", 1 => x"9e", 2 => x"ca", 3 => x"f3"),   -- a89ecaf3
         3 => (0 => x"24", 1 => x"66", 2 => x"ef", 3 => x"97"))   -- 2466ef97
        ),
      1 =>
      (
        0 =>
        -- ae2d8a571e03ac9c9eb76fac45af8e51
        (0 => (0 => x"ae", 1 => x"2d", 2 => x"8a", 3 => x"57"),   -- ae2d8a57
         1 => (0 => x"1e", 1 => x"03", 2 => x"ac", 3 => x"9c"),   -- 1e03ac9c
         2 => (0 => x"9e", 1 => x"b7", 2 => x"6f", 3 => x"ac"),   -- 9eb76fac
         3 => (0 => x"45", 1 => x"af", 2 => x"8e", 3 => x"51")),  -- 45af8e51
        1 =>
        -- f5d3d58503b9699de785895a96fdbaaf
        (0 => (0 => x"f5", 1 => x"d3", 2 => x"d5", 3 => x"85"),   -- f5d3d585
         1 => (0 => x"03", 1 => x"b9", 2 => x"69", 3 => x"9d"),   -- 03b9699d
         2 => (0 => x"e7", 1 => x"85", 2 => x"89", 3 => x"5a"),   -- e785895a
         3 => (0 => x"96", 1 => x"fd", 2 => x"ba", 3 => x"af"))   -- 96fdbaaf
        ),
      2 =>
      (
        0 =>
        -- 30c81c46a35ce411e5fbc1191a0a52ef
        (0 => (0 => x"30", 1 => x"c8", 2 => x"1c", 3 => x"46"),   -- 30c81c46
         1 => (0 => x"a3", 1 => x"5c", 2 => x"e4", 3 => x"11"),   -- a35ce411
         2 => (0 => x"e5", 1 => x"fb", 2 => x"c1", 3 => x"19"),   -- e5fbc119
         3 => (0 => x"1a", 1 => x"0a", 2 => x"52", 3 => x"ef")),  -- 1a0a52ef
        1 =>
        -- 43b1cd7f598ece23881b00e3ed030688
        (0 => (0 => x"43", 1 => x"b1", 2 => x"cd", 3 => x"7f"),   -- 43b1cd7f
         1 => (0 => x"59", 1 => x"8e", 2 => x"ce", 3 => x"23"),   -- 598ece23
         2 => (0 => x"88", 1 => x"1b", 2 => x"00", 3 => x"e3"),   -- 881b00e3
         3 => (0 => x"ed", 1 => x"03", 2 => x"06", 3 => x"88"))   -- ed030688
        ),
      3 =>
      (
        0 =>
        -- f69f2445df4f9b17ad2b417be66c3710
        (0 => (0 => x"f6", 1 => x"9f", 2 => x"24", 3 => x"45"),   -- f69f2445
         1 => (0 => x"df", 1 => x"4f", 2 => x"9b", 3 => x"17"),   -- df4f9b17
         2 => (0 => x"ad", 1 => x"2b", 2 => x"41", 3 => x"7b"),   -- ad2b417b
         3 => (0 => x"e6", 1 => x"6c", 2 => x"37", 3 => x"10")),  -- e66c3710
        1 =>
        -- 7b0c785e27e8ad3f8223207104725dd4
        (0 => (0 => x"7b", 1 => x"0c", 2 => x"78", 3 => x"5e"),   -- 7b0c785e
         1 => (0 => x"27", 1 => x"e8", 2 => x"ad", 3 => x"3f"),   -- 27e8ad3f
         2 => (0 => x"82", 1 => x"23", 2 => x"20", 3 => x"71"),   -- 82232071
         3 => (0 => x"04", 1 => x"72", 2 => x"5d", 3 => x"d4"))   -- 04725dd4
        )
      );


  constant TestVector128_CBC : TestVectorType(0 to 3, 0 to 1)(0 to 4-1)(0 to 4-1)(7 downto 0) :=
    (
      0 =>
      (
        0 =>
        -- 6bc1bee22e409f96e93d7e117393172a
        (0 => (0 => x"6b", 1 => x"c1", 2 => x"be", 3 => x"e2"),   -- 6bc1bee2
         1 => (0 => x"2e", 1 => x"40", 2 => x"9f", 3 => x"96"),   -- 2e409f96
         2 => (0 => x"e9", 1 => x"3d", 2 => x"7e", 3 => x"11"),   -- e93d7e11
         3 => (0 => x"73", 1 => x"93", 2 => x"17", 3 => x"2a")),  -- 7393172a
        1 =>
        -- 7649abac8119b246cee98e9b12e9197d
        (0 => (0 => x"76", 1 => x"49", 2 => x"ab", 3 => x"ac"),   -- 7649abac
         1 => (0 => x"81", 1 => x"19", 2 => x"b2", 3 => x"46"),   -- 8119b246
         2 => (0 => x"ce", 1 => x"e9", 2 => x"8e", 3 => x"9b"),   -- cee98e9b
         3 => (0 => x"12", 1 => x"e9", 2 => x"19", 3 => x"7d"))   -- 12e9197d
        ),
      1 =>
      (
        0 =>
        -- ae2d8a571e03ac9c9eb76fac45af8e51
        (0 => (0 => x"ae", 1 => x"2d", 2 => x"8a", 3 => x"57"),   -- ae2d8a57
         1 => (0 => x"1e", 1 => x"03", 2 => x"ac", 3 => x"9c"),   -- 1e03ac9c
         2 => (0 => x"9e", 1 => x"b7", 2 => x"6f", 3 => x"ac"),   -- 9eb76fac
         3 => (0 => x"45", 1 => x"af", 2 => x"8e", 3 => x"51")),  -- 45af8e51
        1 =>
        -- 5086cb9b507219ee95db113a917678b2
        (0 => (0 => x"50", 1 => x"86", 2 => x"cb", 3 => x"9b"),   -- 5086cb9b
         1 => (0 => x"50", 1 => x"72", 2 => x"19", 3 => x"ee"),   -- 507219ee
         2 => (0 => x"95", 1 => x"db", 2 => x"11", 3 => x"3a"),   -- 95db113a
         3 => (0 => x"91", 1 => x"76", 2 => x"78", 3 => x"b2"))   -- 917678b2
        ),
      2 =>
      (
        0 =>
        -- 30c81c46a35ce411e5fbc1191a0a52ef
        (0 => (0 => x"30", 1 => x"c8", 2 => x"1c", 3 => x"46"),   -- 30c81c46
         1 => (0 => x"a3", 1 => x"5c", 2 => x"e4", 3 => x"11"),   -- a35ce411
         2 => (0 => x"e5", 1 => x"fb", 2 => x"c1", 3 => x"19"),   -- e5fbc119
         3 => (0 => x"1a", 1 => x"0a", 2 => x"52", 3 => x"ef")),  -- 1a0a52ef
        1 =>
        -- 73bed6b8e3c1743b7116e69e22229516
        (0 => (0 => x"73", 1 => x"be", 2 => x"d6", 3 => x"b8"),   -- 73bed6b8
         1 => (0 => x"e3", 1 => x"c1", 2 => x"74", 3 => x"3b"),   -- e3c1743b
         2 => (0 => x"71", 1 => x"16", 2 => x"e6", 3 => x"9e"),   -- 7116e69e
         3 => (0 => x"22", 1 => x"22", 2 => x"95", 3 => x"16"))   -- 22229516
        ),
      3 =>
      (
        0 =>
        -- f69f2445df4f9b17ad2b417be66c3710
        (0 => (0 => x"f6", 1 => x"9f", 2 => x"24", 3 => x"45"),   -- f69f2445
         1 => (0 => x"df", 1 => x"4f", 2 => x"9b", 3 => x"17"),   -- df4f9b17
         2 => (0 => x"ad", 1 => x"2b", 2 => x"41", 3 => x"7b"),   -- ad2b417b
         3 => (0 => x"e6", 1 => x"6c", 2 => x"37", 3 => x"10")),  -- e66c3710
        1 =>
        -- 3ff1caa1681fac09120eca307586e1a7
        (0 => (0 => x"3f", 1 => x"f1", 2 => x"ca", 3 => x"a1"),   -- 3ff1caa1
         1 => (0 => x"68", 1 => x"1f", 2 => x"ac", 3 => x"09"),   -- 681fac09
         2 => (0 => x"12", 1 => x"0e", 2 => x"ca", 3 => x"30"),   -- 120eca30
         3 => (0 => x"75", 1 => x"86", 2 => x"e1", 3 => x"a7"))   -- 7586e1a7
        )
      );


  constant TestVector128_CFB128 : TestVectorType(0 to 3, 0 to 1)(0 to 4-1)(0 to 4-1)(7 downto 0) :=
    (
      0 =>
      (
        0 =>
        -- 6bc1bee22e409f96e93d7e117393172a
        (0 => (0 => x"6b", 1 => x"c1", 2 => x"be", 3 => x"e2"),   -- 6bc1bee2
         1 => (0 => x"2e", 1 => x"40", 2 => x"9f", 3 => x"96"),   -- 2e409f96
         2 => (0 => x"e9", 1 => x"3d", 2 => x"7e", 3 => x"11"),   -- e93d7e11
         3 => (0 => x"73", 1 => x"93", 2 => x"17", 3 => x"2a")),  -- 7393172a
        1 =>
        -- 3b3fd92eb72dad20333449f8e83cfb4a
        (0 => (0 => x"3b", 1 => x"3f", 2 => x"d9", 3 => x"2e"),   -- 3b3fd92e
         1 => (0 => x"b7", 1 => x"2d", 2 => x"ad", 3 => x"20"),   -- b72dad20
         2 => (0 => x"33", 1 => x"34", 2 => x"49", 3 => x"f8"),   -- 333449f8
         3 => (0 => x"e8", 1 => x"3c", 2 => x"fb", 3 => x"4a"))   -- e83cfb4a
        ),
      1 =>
      (
        0 =>
        -- ae2d8a571e03ac9c9eb76fac45af8e51
        (0 => (0 => x"ae", 1 => x"2d", 2 => x"8a", 3 => x"57"),   -- ae2d8a57
         1 => (0 => x"1e", 1 => x"03", 2 => x"ac", 3 => x"9c"),   -- 1e03ac9c
         2 => (0 => x"9e", 1 => x"b7", 2 => x"6f", 3 => x"ac"),   -- 9eb76fac
         3 => (0 => x"45", 1 => x"af", 2 => x"8e", 3 => x"51")),  -- 45af8e51
        1 =>
        -- c8a64537a0b3a93fcde3cdad9f1ce58b
        (0 => (0 => x"c8", 1 => x"a6", 2 => x"45", 3 => x"37"),   -- c8a64537
         1 => (0 => x"a0", 1 => x"b3", 2 => x"a9", 3 => x"3f"),   -- a0b3a93f
         2 => (0 => x"cd", 1 => x"e3", 2 => x"cd", 3 => x"ad"),   -- cde3cdad
         3 => (0 => x"9f", 1 => x"1c", 2 => x"e5", 3 => x"8b"))   -- 9f1ce58b
        ),
      2 =>
      (
        0 =>
        -- 30c81c46a35ce411e5fbc1191a0a52ef
        (0 => (0 => x"30", 1 => x"c8", 2 => x"1c", 3 => x"46"),   -- 30c81c46
         1 => (0 => x"a3", 1 => x"5c", 2 => x"e4", 3 => x"11"),   -- a35ce411
         2 => (0 => x"e5", 1 => x"fb", 2 => x"c1", 3 => x"19"),   -- e5fbc119
         3 => (0 => x"1a", 1 => x"0a", 2 => x"52", 3 => x"ef")),  -- 1a0a52ef
        1 =>
        -- 26751f67a3cbb140b1808cf187a4f4df
        (0 => (0 => x"26", 1 => x"75", 2 => x"1f", 3 => x"67"),   -- 26751f67
         1 => (0 => x"a3", 1 => x"cb", 2 => x"b1", 3 => x"40"),   -- a3cbb140
         2 => (0 => x"b1", 1 => x"80", 2 => x"8c", 3 => x"f1"),   -- b1808cf1
         3 => (0 => x"87", 1 => x"a4", 2 => x"f4", 3 => x"df"))   -- 87a4f4df
        ),
      3 =>
      (
        0 =>
        -- f69f2445df4f9b17ad2b417be66c3710
        (0 => (0 => x"f6", 1 => x"9f", 2 => x"24", 3 => x"45"),   -- f69f2445
         1 => (0 => x"df", 1 => x"4f", 2 => x"9b", 3 => x"17"),   -- df4f9b17
         2 => (0 => x"ad", 1 => x"2b", 2 => x"41", 3 => x"7b"),   -- ad2b417b
         3 => (0 => x"e6", 1 => x"6c", 2 => x"37", 3 => x"10")),  -- e66c3710
        1 =>
        -- c04b05357c5d1c0eeac4c66f9ff7f2e6
        (0 => (0 => x"c0", 1 => x"4b", 2 => x"05", 3 => x"35"),   -- c04b0535
         1 => (0 => x"7c", 1 => x"5d", 2 => x"1c", 3 => x"0e"),   -- 7c5d1c0e
         2 => (0 => x"ea", 1 => x"c4", 2 => x"c6", 3 => x"6f"),   -- eac4c66f
         3 => (0 => x"9f", 1 => x"f7", 2 => x"f2", 3 => x"e6"))   -- 9ff7f2e6
        )
      );


  constant TestVector128_OFB : TestVectorType(0 to 3, 0 to 1)(0 to 4-1)(0 to 4-1)(7 downto 0) :=
    (
      0 =>
      (
        0 =>
        -- 6bc1bee22e409f96e93d7e117393172a
        (0 => (0 => x"6b", 1 => x"c1", 2 => x"be", 3 => x"e2"),   -- 6bc1bee2
         1 => (0 => x"2e", 1 => x"40", 2 => x"9f", 3 => x"96"),   -- 2e409f96
         2 => (0 => x"e9", 1 => x"3d", 2 => x"7e", 3 => x"11"),   -- e93d7e11
         3 => (0 => x"73", 1 => x"93", 2 => x"17", 3 => x"2a")),  -- 7393172a
        1 =>
        -- 3b3fd92eb72dad20333449f8e83cfb4a
        (0 => (0 => x"3b", 1 => x"3f", 2 => x"d9", 3 => x"2e"),   -- 3b3fd92e
         1 => (0 => x"b7", 1 => x"2d", 2 => x"ad", 3 => x"20"),   -- b72dad20
         2 => (0 => x"33", 1 => x"34", 2 => x"49", 3 => x"f8"),   -- 333449f8
         3 => (0 => x"e8", 1 => x"3c", 2 => x"fb", 3 => x"4a"))   -- e83cfb4a
        ),
      1 =>
      (
        0 =>
        -- ae2d8a571e03ac9c9eb76fac45af8e51
        (0 => (0 => x"ae", 1 => x"2d", 2 => x"8a", 3 => x"57"),   -- ae2d8a57
         1 => (0 => x"1e", 1 => x"03", 2 => x"ac", 3 => x"9c"),   -- 1e03ac9c
         2 => (0 => x"9e", 1 => x"b7", 2 => x"6f", 3 => x"ac"),   -- 9eb76fac
         3 => (0 => x"45", 1 => x"af", 2 => x"8e", 3 => x"51")),  -- 45af8e51
        1 =>
        -- 7789508d16918f03f53c52dac54ed825
        (0 => (0 => x"77", 1 => x"89", 2 => x"50", 3 => x"8d"),   -- 7789508d
         1 => (0 => x"16", 1 => x"91", 2 => x"8f", 3 => x"03"),   -- 16918f03
         2 => (0 => x"f5", 1 => x"3c", 2 => x"52", 3 => x"da"),   -- f53c52da
         3 => (0 => x"c5", 1 => x"4e", 2 => x"d8", 3 => x"25"))   -- c54ed825
        ),
      2 =>
      (
        0 =>
        -- 30c81c46a35ce411e5fbc1191a0a52ef
        (0 => (0 => x"30", 1 => x"c8", 2 => x"1c", 3 => x"46"),   -- 30c81c46
         1 => (0 => x"a3", 1 => x"5c", 2 => x"e4", 3 => x"11"),   -- a35ce411
         2 => (0 => x"e5", 1 => x"fb", 2 => x"c1", 3 => x"19"),   -- e5fbc119
         3 => (0 => x"1a", 1 => x"0a", 2 => x"52", 3 => x"ef")),  -- 1a0a52ef
        1 =>
        -- 9740051e9c5fecf64344f7a82260edcc
        (0 => (0 => x"97", 1 => x"40", 2 => x"05", 3 => x"1e"),   -- 9740051e
         1 => (0 => x"9c", 1 => x"5f", 2 => x"ec", 3 => x"f6"),   -- 9c5fecf6
         2 => (0 => x"43", 1 => x"44", 2 => x"f7", 3 => x"a8"),   -- 4344f7a8
         3 => (0 => x"22", 1 => x"60", 2 => x"ed", 3 => x"cc"))   -- 2260edcc
        ),
      3 =>
      (
        0 =>
        -- f69f2445df4f9b17ad2b417be66c3710
        (0 => (0 => x"f6", 1 => x"9f", 2 => x"24", 3 => x"45"),   -- f69f2445
         1 => (0 => x"df", 1 => x"4f", 2 => x"9b", 3 => x"17"),   -- df4f9b17
         2 => (0 => x"ad", 1 => x"2b", 2 => x"41", 3 => x"7b"),   -- ad2b417b
         3 => (0 => x"e6", 1 => x"6c", 2 => x"37", 3 => x"10")),  -- e66c3710
        1 =>
        -- 304c6528f659c77866a510d9c1d6ae5e
        (0 => (0 => x"30", 1 => x"4c", 2 => x"65", 3 => x"28"),   -- 304c6528
         1 => (0 => x"f6", 1 => x"59", 2 => x"c7", 3 => x"78"),   -- f659c778
         2 => (0 => x"66", 1 => x"a5", 2 => x"10", 3 => x"d9"),   -- 66a510d9
         3 => (0 => x"c1", 1 => x"d6", 2 => x"ae", 3 => x"5e"))   -- c1d6ae5e
        )
      );


  constant TestVector128_CTR : TestVectorType(0 to 3, 0 to 1)(0 to 4-1)(0 to 4-1)(7 downto 0) :=
    (
      0 =>
      (
        0 =>
        -- 6bc1bee22e409f96e93d7e117393172a
        (0 => (0 => x"6b", 1 => x"c1", 2 => x"be", 3 => x"e2"),   -- 6bc1bee2
         1 => (0 => x"2e", 1 => x"40", 2 => x"9f", 3 => x"96"),   -- 2e409f96
         2 => (0 => x"e9", 1 => x"3d", 2 => x"7e", 3 => x"11"),   -- e93d7e11
         3 => (0 => x"73", 1 => x"93", 2 => x"17", 3 => x"2a")),  -- 7393172a
        1 =>
        -- 874d6191b620e3261bef6864990db6ce
        (0 => (0 => x"87", 1 => x"4d", 2 => x"61", 3 => x"91"),   -- 874d6191
         1 => (0 => x"b6", 1 => x"20", 2 => x"e3", 3 => x"26"),   -- b620e326
         2 => (0 => x"1b", 1 => x"ef", 2 => x"68", 3 => x"64"),   -- 1bef6864
         3 => (0 => x"99", 1 => x"0d", 2 => x"b6", 3 => x"ce"))   -- 990db6ce
        ),
      1 =>
      (
        0 =>
        -- ae2d8a571e03ac9c9eb76fac45af8e51
        (0 => (0 => x"ae", 1 => x"2d", 2 => x"8a", 3 => x"57"),   -- ae2d8a57
         1 => (0 => x"1e", 1 => x"03", 2 => x"ac", 3 => x"9c"),   -- 1e03ac9c
         2 => (0 => x"9e", 1 => x"b7", 2 => x"6f", 3 => x"ac"),   -- 9eb76fac
         3 => (0 => x"45", 1 => x"af", 2 => x"8e", 3 => x"51")),  -- 45af8e51
        1 =>
        -- 9806f66b7970fdff8617187bb9fffdff
        (0 => (0 => x"98", 1 => x"06", 2 => x"f6", 3 => x"6b"),   -- 9806f66b
         1 => (0 => x"79", 1 => x"70", 2 => x"fd", 3 => x"ff"),   -- 7970fdff
         2 => (0 => x"86", 1 => x"17", 2 => x"18", 3 => x"7b"),   -- 8617187b
         3 => (0 => x"b9", 1 => x"ff", 2 => x"fd", 3 => x"ff"))   -- b9fffdff
        ),
      2 =>
      (
        0 =>
        -- 30c81c46a35ce411e5fbc1191a0a52ef
        (0 => (0 => x"30", 1 => x"c8", 2 => x"1c", 3 => x"46"),   -- 30c81c46
         1 => (0 => x"a3", 1 => x"5c", 2 => x"e4", 3 => x"11"),   -- a35ce411
         2 => (0 => x"e5", 1 => x"fb", 2 => x"c1", 3 => x"19"),   -- e5fbc119
         3 => (0 => x"1a", 1 => x"0a", 2 => x"52", 3 => x"ef")),  -- 1a0a52ef
        1 =>
        -- 5ae4df3edbd5d35e5b4f09020db03eab
        (0 => (0 => x"5a", 1 => x"e4", 2 => x"df", 3 => x"3e"),   -- 5ae4df3e
         1 => (0 => x"db", 1 => x"d5", 2 => x"d3", 3 => x"5e"),   -- dbd5d35e
         2 => (0 => x"5b", 1 => x"4f", 2 => x"09", 3 => x"02"),   -- 5b4f0902
         3 => (0 => x"0d", 1 => x"b0", 2 => x"3e", 3 => x"ab"))   -- 0db03eab
        ),
      3 =>
      (
        0 =>
        -- f69f2445df4f9b17ad2b417be66c3710
        (0 => (0 => x"f6", 1 => x"9f", 2 => x"24", 3 => x"45"),   -- f69f2445
         1 => (0 => x"df", 1 => x"4f", 2 => x"9b", 3 => x"17"),   -- df4f9b17
         2 => (0 => x"ad", 1 => x"2b", 2 => x"41", 3 => x"7b"),   -- ad2b417b
         3 => (0 => x"e6", 1 => x"6c", 2 => x"37", 3 => x"10")),  -- e66c3710
        1 =>
        -- 1e031dda2fbe03d1792170a0f3009cee
        (0 => (0 => x"1e", 1 => x"03", 2 => x"1d", 3 => x"da"),   -- 1e031dda
         1 => (0 => x"2f", 1 => x"be", 2 => x"03", 3 => x"d1"),   -- 2fbe03d1
         2 => (0 => x"79", 1 => x"21", 2 => x"70", 3 => x"a0"),   -- 792170a0
         3 => (0 => x"f3", 1 => x"00", 2 => x"9c", 3 => x"ee"))   -- f3009cee
        )
      );


  constant Sbox    : SboxType(0 to WordRange-1)(Word'range) := InitSbox(WordSize);
  constant InvSbox : SboxType(0 to WordRange-1)(Word'range) := InitInvSbox(Sbox);


begin

  -----------------------------------------------------------------------------
  -- Modes of Operation of the AES taken from:
  -- NIST Special Publication 800-38A Recommendation for Block 2001 Edition
  -- Cipher Modes of Operation, Methods and Techniques
  -----------------------------------------------------------------------------

  process is
    variable State0      : StateType(0 to 4-1)(0 to 4-1)(7 downto 0);
    variable KeySchedule : KeyScheduleType(0 to 15-1)(0 to 4-1)(0 to 4-1)(7 downto 0);
  begin  -- process
    KeySchedule := KeyExpand(Key256, KeySchedule);
    for i in TestVector256_ECB'range loop
      State0 := Encrypt(Sbox, KeySchedule, TestVector256_ECB(i, 0));
      assert State0 = TestVector256_ECB(i, 1)
        report "AES-256 ECB Encrypt failed !!!"
        severity failure;
      State0 := Decrypt(InvSbox, KeySchedule, TestVector256_ECB(i, 1));
      assert State0 = TestVector256_ECB(i, 0)
        report "AES-256 ECB Decrypt failed !!!"
        severity failure;
    end loop;  -- i
    report "AES-256 ECB Encrypt / Decrypt passed.";
    wait;
  end process;

  process is
    variable State0      : StateType(0 to 4-1)(0 to 4-1)(7 downto 0);
    variable KeySchedule : KeyScheduleType(0 to 13-1)(0 to 4-1)(0 to 4-1)(7 downto 0);
  begin  -- process
    KeySchedule := KeyExpand(Key192, KeySchedule);
    for i in TestVector192_ECB'range loop
      State0 := Encrypt(Sbox, KeySchedule, TestVector192_ECB(i, 0));
      assert State0 = TestVector192_ECB(i, 1)
        report "AES-192 ECB Encrypt failed !!!"
        severity failure;
      State0 := Decrypt(InvSbox, KeySchedule, TestVector192_ECB(i, 1));
      assert State0 = TestVector192_ECB(i, 0)
        report "AES-192 ECB Decrypt failed !!!"
        severity failure;
    end loop;  -- i
    report "AES-192 ECB Encrypt / Decrypt passed.";
    wait;
  end process;

  process is
    variable State0      : StateType(0 to 4-1)(0 to 4-1)(7 downto 0);
    variable KeySchedule : KeyScheduleType(0 to 11-1)(0 to 4-1)(0 to 4-1)(7 downto 0);
  begin  -- process
    KeySchedule := KeyExpand(Key128, KeySchedule);
    for i in TestVector128_ECB'range loop
      State0 := Encrypt(Sbox, KeySchedule, TestVector128_ECB(i, 0));
      assert State0 = TestVector128_ECB(i, 1)
        report "AES-128 ECB Encrypt failed !!!"
        severity failure;
      State0 := Decrypt(InvSbox, KeySchedule, TestVector128_ECB(i, 1));
      assert State0 = TestVector128_ECB(i, 0)
        report "AES-128 ECB Decrypt failed !!!"
        severity failure;
    end loop;  -- i
    report "AES-128 ECB Encrypt / Decrypt passed.";
    wait;
  end process;

  process is
    variable State0      : StateType(0 to 4-1)(0 to 4-1)(7 downto 0);
    variable KeySchedule : KeyScheduleType(0 to 15-1)(0 to 4-1)(0 to 4-1)(7 downto 0);
  begin  -- process
    KeySchedule := KeyExpand(Key256, KeySchedule);
    State0      := InitializationVector;
    for i in TestVector256_CBC'range loop
      State0 := Encrypt(Sbox, KeySchedule, TestVector256_CBC(i, 0) + State0);
      assert State0 = TestVector256_CBC(i, 1)
        report "AES-256 CBC Encrypt failed !!!"
        severity failure;
    end loop;  -- i
    State0 := InitializationVector;
    for i in TestVector256_CBC'range loop
      assert Decrypt(InvSbox, KeySchedule, TestVector256_CBC(i, 1)) + State0 = TestVector256_CBC(i, 0)
        report "AES-256 CBC Decrypt failed !!!"
        severity failure;
      State0 := TestVector256_CBC(i, 1);
    end loop;  -- i
    report "AES-256 CBC Encrypt / Decrypt passed.";
    wait;
  end process;

  process is
    variable State0      : StateType(0 to 4-1)(0 to 4-1)(7 downto 0);
    variable KeySchedule : KeyScheduleType(0 to 13-1)(0 to 4-1)(0 to 4-1)(7 downto 0);
  begin  -- process
    KeySchedule := KeyExpand(Key192, KeySchedule);
    State0      := InitializationVector;
    for i in TestVector192_CBC'range loop
      State0 := Encrypt(Sbox, KeySchedule, TestVector192_CBC(i, 0) + State0);
      assert State0 = TestVector192_CBC(i, 1)
        report "AES-192 CBC Encrypt failed !!!"
        severity note;
    end loop;  -- i
    State0 := InitializationVector;
    for i in TestVector192_CBC'range loop
      assert Decrypt(InvSbox, KeySchedule, TestVector192_CBC(i, 1)) + State0 = TestVector192_CBC(i, 0)
        report "AES-192 CBC Decrypt failed !!!"
        severity note;
      State0 := TestVector192_CBC(i, 1);
    end loop;  -- i
    report "AES-192 CBC Encrypt / Decrypt passed.";
    wait;
  end process;

  process is
    variable State0      : StateType(0 to 4-1)(0 to 4-1)(7 downto 0);
    variable KeySchedule : KeyScheduleType(0 to 11-1)(0 to 4-1)(0 to 4-1)(7 downto 0);
  begin  -- process
    KeySchedule := KeyExpand(Key128, KeySchedule);
    State0      := InitializationVector;
    for i in TestVector128_CBC'range loop
      State0 := Encrypt(Sbox, KeySchedule, TestVector128_CBC(i, 0) + State0);
      assert State0 = TestVector128_CBC(i, 1)
        report "AES-128 CBC Encrypt failed !!!"
        severity failure;
    end loop;  -- i
    State0 := InitializationVector;
    for i in TestVector128_CBC'range loop
      assert Decrypt(InvSbox, KeySchedule, TestVector128_CBC(i, 1)) + State0 = TestVector128_CBC(i, 0)
        report "AES-128 CBC Decrypt failed !!!"
        severity failure;
      State0 := TestVector128_CBC(i, 1);
    end loop;  -- i
    report "AES-128 CBC Encrypt / Decrypt passed.";
    wait;
  end process;

  process is
    variable State0      : StateType(0 to 4-1)(0 to 4-1)(7 downto 0);
    variable KeySchedule : KeyScheduleType(0 to 15-1)(0 to 4-1)(0 to 4-1)(7 downto 0);
  begin  -- process
    KeySchedule := KeyExpand(Key256, KeySchedule);
    State0      := InitializationVector;
    for i in TestVector256_CFB128'range loop
      State0 := Encrypt(Sbox, KeySchedule, State0) + TestVector256_CFB128(i, 0);
      assert State0 = TestVector256_CFB128(i, 1)
        report "AES-256 CFB128 Encrypt failed !!!"
        severity failure;
    end loop;  -- i
    State0 := InitializationVector;
    for i in TestVector256_CFB128'range loop
      assert Encrypt(Sbox, KeySchedule, State0) + TestVector256_CFB128(i, 1) = TestVector256_CFB128(i, 0)
        report "AES-256 CFB128 Decrypt failed !!!"
        severity failure;
      State0 := TestVector256_CFB128(i, 1);
    end loop;  -- i
    report "AES-256 CFB128 Encrypt / Decrypt passed.";
    wait;
  end process;

  process is
    variable State0      : StateType(0 to 4-1)(0 to 4-1)(7 downto 0);
    variable KeySchedule : KeyScheduleType(0 to 13-1)(0 to 4-1)(0 to 4-1)(7 downto 0);
  begin  -- process
    KeySchedule := KeyExpand(Key192, KeySchedule);
    State0      := InitializationVector;
    for i in TestVector192_CFB128'range loop
      State0 := Encrypt(Sbox, KeySchedule, State0) + TestVector192_CFB128(i, 0);
      assert State0 = TestVector192_CFB128(i, 1)
        report "AES-192 CFB128 Encrypt failed !!!"
        severity failure;
    end loop;  -- i
    State0 := InitializationVector;
    for i in TestVector192_CFB128'range loop
      assert Encrypt(Sbox, KeySchedule, State0) + TestVector192_CFB128(i, 1) = TestVector192_CFB128(i, 0)
        report "AES-192 CFB128 Decrypt failed !!!"
        severity failure;
      State0 := TestVector192_CFB128(i, 1);
    end loop;  -- i
    report "AES-192 CFB128 Encrypt / Decrypt passed.";
    wait;
  end process;

  process is
    variable State0      : StateType(0 to 4-1)(0 to 4-1)(7 downto 0);
    variable KeySchedule : KeyScheduleType(0 to 11-1)(0 to 4-1)(0 to 4-1)(7 downto 0);
  begin  -- process
    KeySchedule := KeyExpand(Key128, KeySchedule);
    State0      := InitializationVector;
    for i in TestVector128_CFB128'range loop
      State0 := Encrypt(Sbox, KeySchedule, State0) + TestVector128_CFB128(i, 0);
      assert State0 = TestVector128_CFB128(i, 1)
        report "AES-128 CFB128 Encrypt failed !!!"
        severity failure;
    end loop;  -- i
    State0 := InitializationVector;
    for i in TestVector128_CFB128'range loop
      assert Encrypt(Sbox, KeySchedule, State0) + TestVector128_CFB128(i, 1) = TestVector128_CFB128(i, 0)
        report "AES-128 CFB128 Decrypt failed !!!"
        severity failure;
      State0 := TestVector128_CFB128(i, 1);
    end loop;  -- i
    report "AES-128 CFB128 Encrypt / Decrypt passed.";
    wait;
  end process;

  process is
    variable State0      : StateType(0 to 4-1)(0 to 4-1)(7 downto 0);
    variable KeySchedule : KeyScheduleType(0 to 15-1)(0 to 4-1)(0 to 4-1)(7 downto 0);
  begin  -- process
    KeySchedule := KeyExpand(Key256, KeySchedule);
    State0      := InitializationVector;
    for i in TestVector256_OFB'range loop
      assert Encrypt(Sbox, KeySchedule, State0) + TestVector256_OFB(i, 0) = TestVector256_OFB(i, 1)
        report "AES-256 OFB Encrypt failed !!!"
        severity failure;
      State0 := Encrypt(Sbox, KeySchedule, State0);
    end loop;  -- i
    State0 := InitializationVector;
    for i in TestVector256_OFB'range loop
      assert Encrypt(Sbox, KeySchedule, State0) + TestVector256_OFB(i, 1) = TestVector256_OFB(i, 0)
        report "AES-256 OFB Decrypt failed !!!"
        severity failure;
      State0 := Encrypt(Sbox, KeySchedule, State0);
    end loop;  -- i
    report "AES-256 OFB Encrypt / Decrypt passed.";
    wait;
  end process;

  process is
    variable State0      : StateType(0 to 4-1)(0 to 4-1)(7 downto 0);
    variable KeySchedule : KeyScheduleType(0 to 13-1)(0 to 4-1)(0 to 4-1)(7 downto 0);
  begin  -- process
    KeySchedule := KeyExpand(Key192, KeySchedule);
    State0      := InitializationVector;
    for i in TestVector192_OFB'range loop
      assert Encrypt(Sbox, KeySchedule, State0) + TestVector192_OFB(i, 0) = TestVector192_OFB(i, 1)
        report "AES-192 OFB Encrypt failed !!!"
        severity failure;
      State0 := Encrypt(Sbox, KeySchedule, State0);
    end loop;  -- i
    State0 := InitializationVector;
    for i in TestVector192_OFB'range loop
      assert Encrypt(Sbox, KeySchedule, State0) + TestVector192_OFB(i, 1) = TestVector192_OFB(i, 0)
        report "AES-192 OFB Decrypt failed !!!"
        severity failure;
      State0 := Encrypt(Sbox, KeySchedule, State0);
    end loop;  -- i
    report "AES-192 OFB Encrypt / Decrypt passed.";
    wait;
  end process;

  process is
    variable State0      : StateType(0 to 4-1)(0 to 4-1)(7 downto 0);
    variable KeySchedule : KeyScheduleType(0 to 11-1)(0 to 4-1)(0 to 4-1)(7 downto 0);
  begin  -- process
    KeySchedule := KeyExpand(Key128, KeySchedule);
    State0      := InitializationVector;
    for i in TestVector128_OFB'range loop
      assert Encrypt(Sbox, KeySchedule, State0) + TestVector128_OFB(i, 0) = TestVector128_OFB(i, 1)
        report "AES-128 OFB Encrypt failed !!!"
        severity failure;
      State0 := Encrypt(Sbox, KeySchedule, State0);
    end loop;  -- i
    State0 := InitializationVector;
    for i in TestVector128_OFB'range loop
      assert Encrypt(Sbox, KeySchedule, State0) + TestVector128_OFB(i, 1) = TestVector128_OFB(i, 0)
        report "AES-128 OFB Decrypt failed !!!"
        severity failure;
      State0 := Encrypt(Sbox, KeySchedule, State0);
    end loop;  -- i
    report "AES-128 OFB Encrypt / Decrypt passed.";
    wait;
  end process;

  process is
    variable State0      : StateType(0 to 4-1)(0 to 4-1)(7 downto 0);
    variable KeySchedule : KeyScheduleType(0 to 15-1)(0 to 4-1)(0 to 4-1)(7 downto 0);
  begin  -- process
    KeySchedule := KeyExpand(Key256, KeySchedule);
    State0      := InitialCounter;
    for i in TestVector256_CTR'range loop
      assert Encrypt(Sbox, KeySchedule, State0) + TestVector256_CTR(i, 0) = TestVector256_CTR(i, 1)
        report "AES-256 CTR Encrypt failed !!!"
        severity failure;
      State0 := State0 + 1;
    end loop;  -- i
    State0 := InitialCounter;
    for i in TestVector256_CTR'range loop
      assert Encrypt(Sbox, KeySchedule, State0) + TestVector256_CTR(i, 1) = TestVector256_CTR(i, 0)
        report "AES-256 CTR Decrypt failed !!!"
        severity failure;
      State0 := State0 + 1;
    end loop;  -- i
    report "AES-256 CTR Encrypt / Decrypt passed.";
    wait;
  end process;

  process is
    variable State0      : StateType(0 to 4-1)(0 to 4-1)(7 downto 0);
    variable KeySchedule : KeyScheduleType(0 to 13-1)(0 to 4-1)(0 to 4-1)(7 downto 0);
  begin  -- process
    KeySchedule := KeyExpand(Key192, KeySchedule);
    State0      := InitialCounter;
    for i in TestVector192_CTR'range loop
      assert Encrypt(Sbox, KeySchedule, State0) + TestVector192_CTR(i, 0) = TestVector192_CTR(i, 1)
        report "AES-192 CTR Encrypt failed !!!"
        severity failure;
      State0 := State0 + 1;
    end loop;  -- i
    State0 := InitialCounter;
    for i in TestVector192_CTR'range loop
      assert Encrypt(Sbox, KeySchedule, State0) + TestVector192_CTR(i, 1) = TestVector192_CTR(i, 0)
        report "AES-192 CTR Decrypt failed !!!"
        severity failure;
      State0 := State0 + 1;
    end loop;  -- i
    report "AES-192 CTR Encrypt / Decrypt passed.";
    wait;
  end process;

  process is
    variable State0      : StateType(0 to 4-1)(0 to 4-1)(7 downto 0);
    variable KeySchedule : KeyScheduleType(0 to 11-1)(0 to 4-1)(0 to 4-1)(7 downto 0);
  begin  -- process
    KeySchedule := KeyExpand(Key128, KeySchedule);
    State0      := InitialCounter;
    for i in TestVector128_CTR'range loop
      assert Encrypt(Sbox, KeySchedule, State0) + TestVector128_CTR(i, 0) = TestVector128_CTR(i, 1)
        report "AES-128 CTR Encrypt failed !!!"
        severity failure;
      State0 := State0 + 1;
    end loop;  -- i
    State0 := InitialCounter;
    for i in TestVector128_CTR'range loop
      assert Encrypt(Sbox, KeySchedule, State0) + TestVector128_CTR(i, 1) = TestVector128_CTR(i, 0)
        report "AES-128 CTR Decrypt failed !!!"
        severity failure;
      State0 := State0 + 1;
    end loop;  -- i
    report "AES-128 CTR Encrypt / Decrypt passed.";
    wait;
  end process;

end architecture behavior;
